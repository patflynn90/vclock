module ascii

const glyph_map = {
	`0`: [
		'█████',
		'█   █',
		'█   █',
		'█   █',
		'█████',
	]
	`1`: [
		'  ██ ',
		'   █ ',
		'   █ ',
		'   █ ',
		' ████',
	]
	`2`: [
		'█████',
		'    █',
		'█████',
		'█    ',
		'█████',
	]
	`3`: [
		'█████',
		'    █',
		'█████',
		'    █',
		'█████',
	]
	`4`: [
		'█   █',
		'█   █',
		'█████',
		'    █',
		'    █',
	]
	`5`: [
		'█████',
		'█    ',
		'█████',
		'    █',
		'█████',
	]
	`6`: [
		'█████',
		'█    ',
		'█████',
		'█   █',
		'█████',
	]
	`7`: [
		'█████',
		'    █',
		'    █',
		'    █',
		'    █',
	]
	`8`: [
		'█████',
		'█   █',
		'█████',
		'█   █',
		'█████',
	]
	`9`: [
		'█████',
		'█   █',
		'█████',
		'    █',
		'█████',
	]
	`:`: [
		'     ',
		'  █  ',
		'     ',
		'  █  ',
		'     ',
	]
	` `: [
		'     ',
		'     ',
		'     ',
		'     ',
		'     ',
	]
	`A`: [
		'█████',
		'█   █',
		'█████',
		'█   █',
		'█   █',
	]
	`P`: [
		'█████',
		'█   █',
		'█████',
		'█    ',
		'█    ',
	]
	`M`: [
		'██ ██',
		'██ ██',
		'█ █ █',
		'█   █',
		'█   █',
	]
}

pub fn render_string(s string) []string {
	mut lines := []string{len: 5, init: ''}

	for ch in s {
		art := glyph_map[ch] or { glyph_map[` `] }
		for i, row in art {
			lines[i] += row + ' '
		}
	}
	return lines
}

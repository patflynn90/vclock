module cli

pub struct Config {
pub:
	color        string
	centered     bool
	show_date    bool
	blink        bool
	show_seconds bool
}

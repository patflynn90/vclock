module ascii

const digit_art = {
	`0`: [
		'█████',
		'█   █',
		'█   █',
		'█   █',
		'█████',
	]
	`1`: [
		'  ██ ',
		'   █ ',
		'   █ ',
		'   █ ',
		' ████',
	]
	`2`: [
		'█████',
		'    █',
		'█████',
		'█    ',
		'█████',
	]
	`3`: [
		'█████',
		'    █',
		'█████',
		'    █',
		'█████',
	]
	`4`: [
		'█   █',
		'█   █',
		'█████',
		'    █',
		'    █',
	]
	`5`: [
		'█████',
		'█    ',
		'█████',
		'    █',
		'█████',
	]
	`6`: [
		'█████',
		'█    ',
		'█████',
		'█   █',
		'█████',
	]
	`7`: [
		'█████',
		'    █',
		'    █',
		'    █',
		'    █',
	]
	`8`: [
		'█████',
		'█   █',
		'█████',
		'█   █',
		'█████',
	]
	`9`: [
		'█████',
		'█   █',
		'█████',
		'    █',
		'█████',
	]
	`:`: [
		'     ',
		'  █  ',
		'     ',
		'  █  ',
		'     ',
	]
	` `: [
		'     ',
		'     ',
		'     ',
		'     ',
		'     ',
	]
}

pub fn render_string(s string) []string {
	mut lines := []string{len: 5, init: ''}

	for ch in s {
		art := digit_art[ch] or { digit_art[` `] }
		for i, row in art {
			lines[i] += row + ' '
		}
	}
	return lines
}
